[aimspice]
[description]
174
Inversor cu tranzistor
R1 IN B 1K
RC OUT EC 1K
Q1 OUT B 0 TRANZISTOR
.Model TRANZISTOR NPN TR=5e-9 TF=8e-9
VIN IN 0 DC 5 PULSE(0 5 0 1e-9 1e-9 1e-7 2e-7)
VEC EC 0 DC 5 
[dc]
1
VIN
0
5
0.1
[tran]
1e-9
6e-7
0
X
0
[ana]
1 1
0
1 1
1 1 -1 6
3
v(in)
v(b)
v(out)
[end]
