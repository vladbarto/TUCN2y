[aimspice]
[description]
232
Inversor cu NMOS
M3 DD GG OUT OUT n_mos1 L=1U W=1U 
.model n_mos1 nmos vto=2.5
M2 OUT IN 0 0 n_mos2 L=1U W=1U
.model n_mos2 nmos vto=2.5
VIN IN 0 DC 5 PULSE(0 5 0 1e-10 1e-10 1e-9 2e-9)
VGG GG 0 DC 5
VDD DD 0 DC 5
C OUT 0.5p
[dc]
1
VIN
0
5
0.1
[tran]
1e-10
6e-9
X
X
0
[ana]
4 1
0
1 1
1 1 0 5
2
v(out)
v(in)
[end]
