[aimspice]
[description]
159
Redresor Dubla Alternanta
D1 1 2 DiodaSi
D2 0 1 DiodaSi
D3 0 3 DiodaSi
D4 3 2 DiodaSi
.Model DiodaSi D tt = 1e-9
R 2 0 100
VIN 1 3 DC 5 SIN(0 10 1k 0 0)
[tran]
1e-9
6e-3
0
0.00001
0
[ana]
4 1
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
[end]
