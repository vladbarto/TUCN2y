[aimspice]
[description]
169
RedresorCuFiltru
D1 1 out DiodaSi
D2 0 1 DiodaSi
D3 0 3 DiodaSi
D4 3 out DiodaSi
.Model DiodaSi D tt = 1e-9
RL out 0 100
C1 out 0 1m
VIN 1 3 DC 5 sin(0 8 50 0 0)
[tran]
1e-9
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -5.49694E-29 8
1
v(out)
[end]
